/*
ESTE EXEMPLO DESCREVE O NÍVEL 
DE ABSTRAÇÃO ESTRUTURAL DO HDL
*/

module or_base(a, b, c);

input a, b;
output c;

or (c, a, b); // EXEMPLO ESTRUTURAL

endmodule
