library verilog;
use verilog.vl_types.all;
entity tb_cronometro is
end tb_cronometro;
